module tb_Ins_Dec ();
	
endmodule