module tb_fsm (
);  
    logic ... 
    fsm dut (); 
endmodule